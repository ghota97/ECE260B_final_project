##
## LEF for PtnCells ;
## created by Innovus v19.17-s077_1 on Sun Mar  6 22:46:48 2022
##

VERSION 5.8 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO fullchip
  CLASS BLOCK ;
  SIZE 538.390000 BY 538.200000 ;
  FOREIGN fullchip 0.000000 0.000000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 0.150000 0.520000 0.250000 ;
    END
  END clk
  PIN mem_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 534.150000 0.520000 534.250000 ;
    END
  END mem_in[127]
  PIN mem_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 530.550000 0.520000 530.650000 ;
    END
  END mem_in[126]
  PIN mem_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 526.750000 0.520000 526.850000 ;
    END
  END mem_in[125]
  PIN mem_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 523.150000 0.520000 523.250000 ;
    END
  END mem_in[124]
  PIN mem_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 519.350000 0.520000 519.450000 ;
    END
  END mem_in[123]
  PIN mem_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 515.750000 0.520000 515.850000 ;
    END
  END mem_in[122]
  PIN mem_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 512.150000 0.520000 512.250000 ;
    END
  END mem_in[121]
  PIN mem_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 508.350000 0.520000 508.450000 ;
    END
  END mem_in[120]
  PIN mem_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 504.750000 0.520000 504.850000 ;
    END
  END mem_in[119]
  PIN mem_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 500.950000 0.520000 501.050000 ;
    END
  END mem_in[118]
  PIN mem_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 497.350000 0.520000 497.450000 ;
    END
  END mem_in[117]
  PIN mem_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 493.550000 0.520000 493.650000 ;
    END
  END mem_in[116]
  PIN mem_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 489.950000 0.520000 490.050000 ;
    END
  END mem_in[115]
  PIN mem_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 486.350000 0.520000 486.450000 ;
    END
  END mem_in[114]
  PIN mem_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 482.550000 0.520000 482.650000 ;
    END
  END mem_in[113]
  PIN mem_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 478.950000 0.520000 479.050000 ;
    END
  END mem_in[112]
  PIN mem_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 475.150000 0.520000 475.250000 ;
    END
  END mem_in[111]
  PIN mem_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 471.550000 0.520000 471.650000 ;
    END
  END mem_in[110]
  PIN mem_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 467.950000 0.520000 468.050000 ;
    END
  END mem_in[109]
  PIN mem_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 464.150000 0.520000 464.250000 ;
    END
  END mem_in[108]
  PIN mem_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 460.550000 0.520000 460.650000 ;
    END
  END mem_in[107]
  PIN mem_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 456.750000 0.520000 456.850000 ;
    END
  END mem_in[106]
  PIN mem_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 453.150000 0.520000 453.250000 ;
    END
  END mem_in[105]
  PIN mem_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 449.350000 0.520000 449.450000 ;
    END
  END mem_in[104]
  PIN mem_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 445.750000 0.520000 445.850000 ;
    END
  END mem_in[103]
  PIN mem_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 442.150000 0.520000 442.250000 ;
    END
  END mem_in[102]
  PIN mem_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 438.350000 0.520000 438.450000 ;
    END
  END mem_in[101]
  PIN mem_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 434.750000 0.520000 434.850000 ;
    END
  END mem_in[100]
  PIN mem_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 430.950000 0.520000 431.050000 ;
    END
  END mem_in[99]
  PIN mem_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 427.350000 0.520000 427.450000 ;
    END
  END mem_in[98]
  PIN mem_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 423.750000 0.520000 423.850000 ;
    END
  END mem_in[97]
  PIN mem_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 419.950000 0.520000 420.050000 ;
    END
  END mem_in[96]
  PIN mem_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 416.350000 0.520000 416.450000 ;
    END
  END mem_in[95]
  PIN mem_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 412.550000 0.520000 412.650000 ;
    END
  END mem_in[94]
  PIN mem_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 408.950000 0.520000 409.050000 ;
    END
  END mem_in[93]
  PIN mem_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 405.150000 0.520000 405.250000 ;
    END
  END mem_in[92]
  PIN mem_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 401.550000 0.520000 401.650000 ;
    END
  END mem_in[91]
  PIN mem_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 397.950000 0.520000 398.050000 ;
    END
  END mem_in[90]
  PIN mem_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 394.150000 0.520000 394.250000 ;
    END
  END mem_in[89]
  PIN mem_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 390.550000 0.520000 390.650000 ;
    END
  END mem_in[88]
  PIN mem_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 386.750000 0.520000 386.850000 ;
    END
  END mem_in[87]
  PIN mem_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 383.150000 0.520000 383.250000 ;
    END
  END mem_in[86]
  PIN mem_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 379.550000 0.520000 379.650000 ;
    END
  END mem_in[85]
  PIN mem_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 375.750000 0.520000 375.850000 ;
    END
  END mem_in[84]
  PIN mem_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 372.150000 0.520000 372.250000 ;
    END
  END mem_in[83]
  PIN mem_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 368.350000 0.520000 368.450000 ;
    END
  END mem_in[82]
  PIN mem_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 364.750000 0.520000 364.850000 ;
    END
  END mem_in[81]
  PIN mem_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 360.950000 0.520000 361.050000 ;
    END
  END mem_in[80]
  PIN mem_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 357.350000 0.520000 357.450000 ;
    END
  END mem_in[79]
  PIN mem_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 353.750000 0.520000 353.850000 ;
    END
  END mem_in[78]
  PIN mem_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 349.950000 0.520000 350.050000 ;
    END
  END mem_in[77]
  PIN mem_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 346.350000 0.520000 346.450000 ;
    END
  END mem_in[76]
  PIN mem_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 342.550000 0.520000 342.650000 ;
    END
  END mem_in[75]
  PIN mem_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 338.950000 0.520000 339.050000 ;
    END
  END mem_in[74]
  PIN mem_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 335.350000 0.520000 335.450000 ;
    END
  END mem_in[73]
  PIN mem_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 331.550000 0.520000 331.650000 ;
    END
  END mem_in[72]
  PIN mem_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 327.950000 0.520000 328.050000 ;
    END
  END mem_in[71]
  PIN mem_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 324.150000 0.520000 324.250000 ;
    END
  END mem_in[70]
  PIN mem_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 320.550000 0.520000 320.650000 ;
    END
  END mem_in[69]
  PIN mem_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 316.750000 0.520000 316.850000 ;
    END
  END mem_in[68]
  PIN mem_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 313.150000 0.520000 313.250000 ;
    END
  END mem_in[67]
  PIN mem_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 309.550000 0.520000 309.650000 ;
    END
  END mem_in[66]
  PIN mem_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 305.750000 0.520000 305.850000 ;
    END
  END mem_in[65]
  PIN mem_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 302.150000 0.520000 302.250000 ;
    END
  END mem_in[64]
  PIN mem_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 298.350000 0.520000 298.450000 ;
    END
  END mem_in[63]
  PIN mem_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 294.750000 0.520000 294.850000 ;
    END
  END mem_in[62]
  PIN mem_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 291.150000 0.520000 291.250000 ;
    END
  END mem_in[61]
  PIN mem_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 287.350000 0.520000 287.450000 ;
    END
  END mem_in[60]
  PIN mem_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 283.750000 0.520000 283.850000 ;
    END
  END mem_in[59]
  PIN mem_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 279.950000 0.520000 280.050000 ;
    END
  END mem_in[58]
  PIN mem_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 276.350000 0.520000 276.450000 ;
    END
  END mem_in[57]
  PIN mem_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 272.550000 0.520000 272.650000 ;
    END
  END mem_in[56]
  PIN mem_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 268.950000 0.520000 269.050000 ;
    END
  END mem_in[55]
  PIN mem_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 265.350000 0.520000 265.450000 ;
    END
  END mem_in[54]
  PIN mem_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 261.550000 0.520000 261.650000 ;
    END
  END mem_in[53]
  PIN mem_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 257.950000 0.520000 258.050000 ;
    END
  END mem_in[52]
  PIN mem_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 254.150000 0.520000 254.250000 ;
    END
  END mem_in[51]
  PIN mem_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 250.550000 0.520000 250.650000 ;
    END
  END mem_in[50]
  PIN mem_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 246.750000 0.520000 246.850000 ;
    END
  END mem_in[49]
  PIN mem_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 243.150000 0.520000 243.250000 ;
    END
  END mem_in[48]
  PIN mem_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 239.550000 0.520000 239.650000 ;
    END
  END mem_in[47]
  PIN mem_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 235.750000 0.520000 235.850000 ;
    END
  END mem_in[46]
  PIN mem_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 232.150000 0.520000 232.250000 ;
    END
  END mem_in[45]
  PIN mem_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 228.350000 0.520000 228.450000 ;
    END
  END mem_in[44]
  PIN mem_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 224.750000 0.520000 224.850000 ;
    END
  END mem_in[43]
  PIN mem_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 221.150000 0.520000 221.250000 ;
    END
  END mem_in[42]
  PIN mem_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 217.350000 0.520000 217.450000 ;
    END
  END mem_in[41]
  PIN mem_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 213.750000 0.520000 213.850000 ;
    END
  END mem_in[40]
  PIN mem_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 209.950000 0.520000 210.050000 ;
    END
  END mem_in[39]
  PIN mem_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 206.350000 0.520000 206.450000 ;
    END
  END mem_in[38]
  PIN mem_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 202.550000 0.520000 202.650000 ;
    END
  END mem_in[37]
  PIN mem_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 198.950000 0.520000 199.050000 ;
    END
  END mem_in[36]
  PIN mem_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 195.350000 0.520000 195.450000 ;
    END
  END mem_in[35]
  PIN mem_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 191.550000 0.520000 191.650000 ;
    END
  END mem_in[34]
  PIN mem_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 187.950000 0.520000 188.050000 ;
    END
  END mem_in[33]
  PIN mem_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 184.150000 0.520000 184.250000 ;
    END
  END mem_in[32]
  PIN mem_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 180.550000 0.520000 180.650000 ;
    END
  END mem_in[31]
  PIN mem_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 176.950000 0.520000 177.050000 ;
    END
  END mem_in[30]
  PIN mem_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 173.150000 0.520000 173.250000 ;
    END
  END mem_in[29]
  PIN mem_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 169.550000 0.520000 169.650000 ;
    END
  END mem_in[28]
  PIN mem_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 165.750000 0.520000 165.850000 ;
    END
  END mem_in[27]
  PIN mem_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 162.150000 0.520000 162.250000 ;
    END
  END mem_in[26]
  PIN mem_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 158.350000 0.520000 158.450000 ;
    END
  END mem_in[25]
  PIN mem_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 154.750000 0.520000 154.850000 ;
    END
  END mem_in[24]
  PIN mem_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 151.150000 0.520000 151.250000 ;
    END
  END mem_in[23]
  PIN mem_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 147.350000 0.520000 147.450000 ;
    END
  END mem_in[22]
  PIN mem_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 143.750000 0.520000 143.850000 ;
    END
  END mem_in[21]
  PIN mem_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 139.950000 0.520000 140.050000 ;
    END
  END mem_in[20]
  PIN mem_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 136.350000 0.520000 136.450000 ;
    END
  END mem_in[19]
  PIN mem_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 132.750000 0.520000 132.850000 ;
    END
  END mem_in[18]
  PIN mem_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 128.950000 0.520000 129.050000 ;
    END
  END mem_in[17]
  PIN mem_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 125.350000 0.520000 125.450000 ;
    END
  END mem_in[16]
  PIN mem_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 121.550000 0.520000 121.650000 ;
    END
  END mem_in[15]
  PIN mem_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 117.950000 0.520000 118.050000 ;
    END
  END mem_in[14]
  PIN mem_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 114.150000 0.520000 114.250000 ;
    END
  END mem_in[13]
  PIN mem_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 110.550000 0.520000 110.650000 ;
    END
  END mem_in[12]
  PIN mem_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 106.950000 0.520000 107.050000 ;
    END
  END mem_in[11]
  PIN mem_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 103.150000 0.520000 103.250000 ;
    END
  END mem_in[10]
  PIN mem_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 99.550000 0.520000 99.650000 ;
    END
  END mem_in[9]
  PIN mem_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 95.750000 0.520000 95.850000 ;
    END
  END mem_in[8]
  PIN mem_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 92.150000 0.520000 92.250000 ;
    END
  END mem_in[7]
  PIN mem_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 88.550000 0.520000 88.650000 ;
    END
  END mem_in[6]
  PIN mem_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 84.750000 0.520000 84.850000 ;
    END
  END mem_in[5]
  PIN mem_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 81.150000 0.520000 81.250000 ;
    END
  END mem_in[4]
  PIN mem_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 77.350000 0.520000 77.450000 ;
    END
  END mem_in[3]
  PIN mem_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 73.750000 0.520000 73.850000 ;
    END
  END mem_in[2]
  PIN mem_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 69.950000 0.520000 70.050000 ;
    END
  END mem_in[1]
  PIN mem_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 66.350000 0.520000 66.450000 ;
    END
  END mem_in[0]
  PIN out[159]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.650000 0.000000 0.750000 0.520000 ;
    END
  END out[159]
  PIN out[158]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 3.450000 0.000000 3.550000 0.520000 ;
    END
  END out[158]
  PIN out[157]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 6.850000 0.000000 6.950000 0.520000 ;
    END
  END out[157]
  PIN out[156]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10.250000 0.000000 10.350000 0.520000 ;
    END
  END out[156]
  PIN out[155]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 13.650000 0.000000 13.750000 0.520000 ;
    END
  END out[155]
  PIN out[154]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 17.050000 0.000000 17.150000 0.520000 ;
    END
  END out[154]
  PIN out[153]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 20.450000 0.000000 20.550000 0.520000 ;
    END
  END out[153]
  PIN out[152]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 23.850000 0.000000 23.950000 0.520000 ;
    END
  END out[152]
  PIN out[151]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 27.250000 0.000000 27.350000 0.520000 ;
    END
  END out[151]
  PIN out[150]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 30.650000 0.000000 30.750000 0.520000 ;
    END
  END out[150]
  PIN out[149]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 34.050000 0.000000 34.150000 0.520000 ;
    END
  END out[149]
  PIN out[148]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 37.450000 0.000000 37.550000 0.520000 ;
    END
  END out[148]
  PIN out[147]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 40.850000 0.000000 40.950000 0.520000 ;
    END
  END out[147]
  PIN out[146]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 44.250000 0.000000 44.350000 0.520000 ;
    END
  END out[146]
  PIN out[145]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 47.450000 0.000000 47.550000 0.520000 ;
    END
  END out[145]
  PIN out[144]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 50.850000 0.000000 50.950000 0.520000 ;
    END
  END out[144]
  PIN out[143]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 54.250000 0.000000 54.350000 0.520000 ;
    END
  END out[143]
  PIN out[142]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 57.650000 0.000000 57.750000 0.520000 ;
    END
  END out[142]
  PIN out[141]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 61.050000 0.000000 61.150000 0.520000 ;
    END
  END out[141]
  PIN out[140]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 64.450000 0.000000 64.550000 0.520000 ;
    END
  END out[140]
  PIN out[139]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 67.850000 0.000000 67.950000 0.520000 ;
    END
  END out[139]
  PIN out[138]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 71.250000 0.000000 71.350000 0.520000 ;
    END
  END out[138]
  PIN out[137]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 74.650000 0.000000 74.750000 0.520000 ;
    END
  END out[137]
  PIN out[136]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 78.050000 0.000000 78.150000 0.520000 ;
    END
  END out[136]
  PIN out[135]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 81.450000 0.000000 81.550000 0.520000 ;
    END
  END out[135]
  PIN out[134]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 84.850000 0.000000 84.950000 0.520000 ;
    END
  END out[134]
  PIN out[133]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 88.250000 0.000000 88.350000 0.520000 ;
    END
  END out[133]
  PIN out[132]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 91.450000 0.000000 91.550000 0.520000 ;
    END
  END out[132]
  PIN out[131]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 94.850000 0.000000 94.950000 0.520000 ;
    END
  END out[131]
  PIN out[130]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 98.250000 0.000000 98.350000 0.520000 ;
    END
  END out[130]
  PIN out[129]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 101.650000 0.000000 101.750000 0.520000 ;
    END
  END out[129]
  PIN out[128]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 105.050000 0.000000 105.150000 0.520000 ;
    END
  END out[128]
  PIN out[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 108.450000 0.000000 108.550000 0.520000 ;
    END
  END out[127]
  PIN out[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 111.850000 0.000000 111.950000 0.520000 ;
    END
  END out[126]
  PIN out[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 115.250000 0.000000 115.350000 0.520000 ;
    END
  END out[125]
  PIN out[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 118.650000 0.000000 118.750000 0.520000 ;
    END
  END out[124]
  PIN out[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 122.050000 0.000000 122.150000 0.520000 ;
    END
  END out[123]
  PIN out[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 125.450000 0.000000 125.550000 0.520000 ;
    END
  END out[122]
  PIN out[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 128.850000 0.000000 128.950000 0.520000 ;
    END
  END out[121]
  PIN out[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 132.250000 0.000000 132.350000 0.520000 ;
    END
  END out[120]
  PIN out[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 135.450000 0.000000 135.550000 0.520000 ;
    END
  END out[119]
  PIN out[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 138.850000 0.000000 138.950000 0.520000 ;
    END
  END out[118]
  PIN out[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 142.250000 0.000000 142.350000 0.520000 ;
    END
  END out[117]
  PIN out[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 145.650000 0.000000 145.750000 0.520000 ;
    END
  END out[116]
  PIN out[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 149.050000 0.000000 149.150000 0.520000 ;
    END
  END out[115]
  PIN out[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 152.450000 0.000000 152.550000 0.520000 ;
    END
  END out[114]
  PIN out[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 155.850000 0.000000 155.950000 0.520000 ;
    END
  END out[113]
  PIN out[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 159.250000 0.000000 159.350000 0.520000 ;
    END
  END out[112]
  PIN out[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 162.650000 0.000000 162.750000 0.520000 ;
    END
  END out[111]
  PIN out[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 166.050000 0.000000 166.150000 0.520000 ;
    END
  END out[110]
  PIN out[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 169.450000 0.000000 169.550000 0.520000 ;
    END
  END out[109]
  PIN out[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 172.850000 0.000000 172.950000 0.520000 ;
    END
  END out[108]
  PIN out[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 176.250000 0.000000 176.350000 0.520000 ;
    END
  END out[107]
  PIN out[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 179.650000 0.000000 179.750000 0.520000 ;
    END
  END out[106]
  PIN out[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 182.850000 0.000000 182.950000 0.520000 ;
    END
  END out[105]
  PIN out[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 186.250000 0.000000 186.350000 0.520000 ;
    END
  END out[104]
  PIN out[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 189.650000 0.000000 189.750000 0.520000 ;
    END
  END out[103]
  PIN out[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 193.050000 0.000000 193.150000 0.520000 ;
    END
  END out[102]
  PIN out[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 196.450000 0.000000 196.550000 0.520000 ;
    END
  END out[101]
  PIN out[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 199.850000 0.000000 199.950000 0.520000 ;
    END
  END out[100]
  PIN out[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 203.250000 0.000000 203.350000 0.520000 ;
    END
  END out[99]
  PIN out[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 206.650000 0.000000 206.750000 0.520000 ;
    END
  END out[98]
  PIN out[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 210.050000 0.000000 210.150000 0.520000 ;
    END
  END out[97]
  PIN out[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 213.450000 0.000000 213.550000 0.520000 ;
    END
  END out[96]
  PIN out[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 216.850000 0.000000 216.950000 0.520000 ;
    END
  END out[95]
  PIN out[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 220.250000 0.000000 220.350000 0.520000 ;
    END
  END out[94]
  PIN out[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 223.650000 0.000000 223.750000 0.520000 ;
    END
  END out[93]
  PIN out[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 226.850000 0.000000 226.950000 0.520000 ;
    END
  END out[92]
  PIN out[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 230.250000 0.000000 230.350000 0.520000 ;
    END
  END out[91]
  PIN out[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 233.650000 0.000000 233.750000 0.520000 ;
    END
  END out[90]
  PIN out[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 237.050000 0.000000 237.150000 0.520000 ;
    END
  END out[89]
  PIN out[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 240.450000 0.000000 240.550000 0.520000 ;
    END
  END out[88]
  PIN out[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 243.850000 0.000000 243.950000 0.520000 ;
    END
  END out[87]
  PIN out[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 247.250000 0.000000 247.350000 0.520000 ;
    END
  END out[86]
  PIN out[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 250.650000 0.000000 250.750000 0.520000 ;
    END
  END out[85]
  PIN out[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 254.050000 0.000000 254.150000 0.520000 ;
    END
  END out[84]
  PIN out[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 257.450000 0.000000 257.550000 0.520000 ;
    END
  END out[83]
  PIN out[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 260.850000 0.000000 260.950000 0.520000 ;
    END
  END out[82]
  PIN out[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 264.250000 0.000000 264.350000 0.520000 ;
    END
  END out[81]
  PIN out[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 267.650000 0.000000 267.750000 0.520000 ;
    END
  END out[80]
  PIN out[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 270.850000 0.000000 270.950000 0.520000 ;
    END
  END out[79]
  PIN out[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 274.250000 0.000000 274.350000 0.520000 ;
    END
  END out[78]
  PIN out[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 277.650000 0.000000 277.750000 0.520000 ;
    END
  END out[77]
  PIN out[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 281.050000 0.000000 281.150000 0.520000 ;
    END
  END out[76]
  PIN out[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 284.450000 0.000000 284.550000 0.520000 ;
    END
  END out[75]
  PIN out[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 287.850000 0.000000 287.950000 0.520000 ;
    END
  END out[74]
  PIN out[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 291.250000 0.000000 291.350000 0.520000 ;
    END
  END out[73]
  PIN out[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 294.650000 0.000000 294.750000 0.520000 ;
    END
  END out[72]
  PIN out[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 298.050000 0.000000 298.150000 0.520000 ;
    END
  END out[71]
  PIN out[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 301.450000 0.000000 301.550000 0.520000 ;
    END
  END out[70]
  PIN out[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 304.850000 0.000000 304.950000 0.520000 ;
    END
  END out[69]
  PIN out[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 308.250000 0.000000 308.350000 0.520000 ;
    END
  END out[68]
  PIN out[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 311.650000 0.000000 311.750000 0.520000 ;
    END
  END out[67]
  PIN out[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 314.850000 0.000000 314.950000 0.520000 ;
    END
  END out[66]
  PIN out[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 318.250000 0.000000 318.350000 0.520000 ;
    END
  END out[65]
  PIN out[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 321.650000 0.000000 321.750000 0.520000 ;
    END
  END out[64]
  PIN out[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 325.050000 0.000000 325.150000 0.520000 ;
    END
  END out[63]
  PIN out[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 328.450000 0.000000 328.550000 0.520000 ;
    END
  END out[62]
  PIN out[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 331.850000 0.000000 331.950000 0.520000 ;
    END
  END out[61]
  PIN out[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 335.250000 0.000000 335.350000 0.520000 ;
    END
  END out[60]
  PIN out[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 338.650000 0.000000 338.750000 0.520000 ;
    END
  END out[59]
  PIN out[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 342.050000 0.000000 342.150000 0.520000 ;
    END
  END out[58]
  PIN out[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 345.450000 0.000000 345.550000 0.520000 ;
    END
  END out[57]
  PIN out[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 348.850000 0.000000 348.950000 0.520000 ;
    END
  END out[56]
  PIN out[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 352.250000 0.000000 352.350000 0.520000 ;
    END
  END out[55]
  PIN out[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 355.650000 0.000000 355.750000 0.520000 ;
    END
  END out[54]
  PIN out[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 359.050000 0.000000 359.150000 0.520000 ;
    END
  END out[53]
  PIN out[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 362.250000 0.000000 362.350000 0.520000 ;
    END
  END out[52]
  PIN out[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 365.650000 0.000000 365.750000 0.520000 ;
    END
  END out[51]
  PIN out[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 369.050000 0.000000 369.150000 0.520000 ;
    END
  END out[50]
  PIN out[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 372.450000 0.000000 372.550000 0.520000 ;
    END
  END out[49]
  PIN out[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 375.850000 0.000000 375.950000 0.520000 ;
    END
  END out[48]
  PIN out[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 379.250000 0.000000 379.350000 0.520000 ;
    END
  END out[47]
  PIN out[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 382.650000 0.000000 382.750000 0.520000 ;
    END
  END out[46]
  PIN out[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 386.050000 0.000000 386.150000 0.520000 ;
    END
  END out[45]
  PIN out[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 389.450000 0.000000 389.550000 0.520000 ;
    END
  END out[44]
  PIN out[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 392.850000 0.000000 392.950000 0.520000 ;
    END
  END out[43]
  PIN out[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 396.250000 0.000000 396.350000 0.520000 ;
    END
  END out[42]
  PIN out[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 399.650000 0.000000 399.750000 0.520000 ;
    END
  END out[41]
  PIN out[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 403.050000 0.000000 403.150000 0.520000 ;
    END
  END out[40]
  PIN out[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 406.250000 0.000000 406.350000 0.520000 ;
    END
  END out[39]
  PIN out[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 409.650000 0.000000 409.750000 0.520000 ;
    END
  END out[38]
  PIN out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 413.050000 0.000000 413.150000 0.520000 ;
    END
  END out[37]
  PIN out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 416.450000 0.000000 416.550000 0.520000 ;
    END
  END out[36]
  PIN out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 419.850000 0.000000 419.950000 0.520000 ;
    END
  END out[35]
  PIN out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 423.250000 0.000000 423.350000 0.520000 ;
    END
  END out[34]
  PIN out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 426.650000 0.000000 426.750000 0.520000 ;
    END
  END out[33]
  PIN out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 430.050000 0.000000 430.150000 0.520000 ;
    END
  END out[32]
  PIN out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 433.450000 0.000000 433.550000 0.520000 ;
    END
  END out[31]
  PIN out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 436.850000 0.000000 436.950000 0.520000 ;
    END
  END out[30]
  PIN out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 440.250000 0.000000 440.350000 0.520000 ;
    END
  END out[29]
  PIN out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 443.650000 0.000000 443.750000 0.520000 ;
    END
  END out[28]
  PIN out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 447.050000 0.000000 447.150000 0.520000 ;
    END
  END out[27]
  PIN out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 450.250000 0.000000 450.350000 0.520000 ;
    END
  END out[26]
  PIN out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 453.650000 0.000000 453.750000 0.520000 ;
    END
  END out[25]
  PIN out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 457.050000 0.000000 457.150000 0.520000 ;
    END
  END out[24]
  PIN out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 460.450000 0.000000 460.550000 0.520000 ;
    END
  END out[23]
  PIN out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 463.850000 0.000000 463.950000 0.520000 ;
    END
  END out[22]
  PIN out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 467.250000 0.000000 467.350000 0.520000 ;
    END
  END out[21]
  PIN out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 470.650000 0.000000 470.750000 0.520000 ;
    END
  END out[20]
  PIN out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 474.050000 0.000000 474.150000 0.520000 ;
    END
  END out[19]
  PIN out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 477.450000 0.000000 477.550000 0.520000 ;
    END
  END out[18]
  PIN out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 480.850000 0.000000 480.950000 0.520000 ;
    END
  END out[17]
  PIN out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 484.250000 0.000000 484.350000 0.520000 ;
    END
  END out[16]
  PIN out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 487.650000 0.000000 487.750000 0.520000 ;
    END
  END out[15]
  PIN out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 491.050000 0.000000 491.150000 0.520000 ;
    END
  END out[14]
  PIN out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 494.250000 0.000000 494.350000 0.520000 ;
    END
  END out[13]
  PIN out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 497.650000 0.000000 497.750000 0.520000 ;
    END
  END out[12]
  PIN out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 501.050000 0.000000 501.150000 0.520000 ;
    END
  END out[11]
  PIN out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 504.450000 0.000000 504.550000 0.520000 ;
    END
  END out[10]
  PIN out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 507.850000 0.000000 507.950000 0.520000 ;
    END
  END out[9]
  PIN out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 511.250000 0.000000 511.350000 0.520000 ;
    END
  END out[8]
  PIN out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 514.650000 0.000000 514.750000 0.520000 ;
    END
  END out[7]
  PIN out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 518.050000 0.000000 518.150000 0.520000 ;
    END
  END out[6]
  PIN out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 521.450000 0.000000 521.550000 0.520000 ;
    END
  END out[5]
  PIN out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 524.850000 0.000000 524.950000 0.520000 ;
    END
  END out[4]
  PIN out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 528.250000 0.000000 528.350000 0.520000 ;
    END
  END out[3]
  PIN out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 531.650000 0.000000 531.750000 0.520000 ;
    END
  END out[2]
  PIN out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 535.050000 0.000000 535.150000 0.520000 ;
    END
  END out[1]
  PIN out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 538.250000 0.000000 538.350000 0.520000 ;
    END
  END out[0]
  PIN inst[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 62.750000 0.520000 62.850000 ;
    END
  END inst[16]
  PIN inst[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 58.950000 0.520000 59.050000 ;
    END
  END inst[15]
  PIN inst[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 55.350000 0.520000 55.450000 ;
    END
  END inst[14]
  PIN inst[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 51.550000 0.520000 51.650000 ;
    END
  END inst[13]
  PIN inst[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 47.950000 0.520000 48.050000 ;
    END
  END inst[12]
  PIN inst[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 44.350000 0.520000 44.450000 ;
    END
  END inst[11]
  PIN inst[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 40.550000 0.520000 40.650000 ;
    END
  END inst[10]
  PIN inst[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 36.950000 0.520000 37.050000 ;
    END
  END inst[9]
  PIN inst[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 33.150000 0.520000 33.250000 ;
    END
  END inst[8]
  PIN inst[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 29.550000 0.520000 29.650000 ;
    END
  END inst[7]
  PIN inst[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 25.750000 0.520000 25.850000 ;
    END
  END inst[6]
  PIN inst[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 22.150000 0.520000 22.250000 ;
    END
  END inst[5]
  PIN inst[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 18.550000 0.520000 18.650000 ;
    END
  END inst[4]
  PIN inst[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 14.750000 0.520000 14.850000 ;
    END
  END inst[3]
  PIN inst[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 11.150000 0.520000 11.250000 ;
    END
  END inst[2]
  PIN inst[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 7.350000 0.520000 7.450000 ;
    END
  END inst[1]
  PIN inst[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 3.750000 0.520000 3.850000 ;
    END
  END inst[0]
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.000000 537.750000 0.520000 537.850000 ;
    END
  END reset
  OBS
    LAYER M1 ;
      RECT 0.000000 0.000000 538.390000 538.200000 ;
    LAYER M2 ;
      RECT 0.000000 0.000000 538.390000 538.200000 ;
    LAYER M3 ;
      RECT 0.000000 0.000000 538.390000 538.200000 ;
    LAYER M4 ;
      RECT 0.000000 538.010000 538.390000 538.200000 ;
      RECT 0.680000 537.590000 538.390000 538.010000 ;
      RECT 0.000000 534.410000 538.390000 537.590000 ;
      RECT 0.680000 533.990000 538.390000 534.410000 ;
      RECT 0.000000 530.810000 538.390000 533.990000 ;
      RECT 0.680000 530.390000 538.390000 530.810000 ;
      RECT 0.000000 527.010000 538.390000 530.390000 ;
      RECT 0.680000 526.590000 538.390000 527.010000 ;
      RECT 0.000000 523.410000 538.390000 526.590000 ;
      RECT 0.680000 522.990000 538.390000 523.410000 ;
      RECT 0.000000 519.610000 538.390000 522.990000 ;
      RECT 0.680000 519.190000 538.390000 519.610000 ;
      RECT 0.000000 516.010000 538.390000 519.190000 ;
      RECT 0.680000 515.590000 538.390000 516.010000 ;
      RECT 0.000000 512.410000 538.390000 515.590000 ;
      RECT 0.680000 511.990000 538.390000 512.410000 ;
      RECT 0.000000 508.610000 538.390000 511.990000 ;
      RECT 0.680000 508.190000 538.390000 508.610000 ;
      RECT 0.000000 505.010000 538.390000 508.190000 ;
      RECT 0.680000 504.590000 538.390000 505.010000 ;
      RECT 0.000000 501.210000 538.390000 504.590000 ;
      RECT 0.680000 500.790000 538.390000 501.210000 ;
      RECT 0.000000 497.610000 538.390000 500.790000 ;
      RECT 0.680000 497.190000 538.390000 497.610000 ;
      RECT 0.000000 493.810000 538.390000 497.190000 ;
      RECT 0.680000 493.390000 538.390000 493.810000 ;
      RECT 0.000000 490.210000 538.390000 493.390000 ;
      RECT 0.680000 489.790000 538.390000 490.210000 ;
      RECT 0.000000 486.610000 538.390000 489.790000 ;
      RECT 0.680000 486.190000 538.390000 486.610000 ;
      RECT 0.000000 482.810000 538.390000 486.190000 ;
      RECT 0.680000 482.390000 538.390000 482.810000 ;
      RECT 0.000000 479.210000 538.390000 482.390000 ;
      RECT 0.680000 478.790000 538.390000 479.210000 ;
      RECT 0.000000 475.410000 538.390000 478.790000 ;
      RECT 0.680000 474.990000 538.390000 475.410000 ;
      RECT 0.000000 471.810000 538.390000 474.990000 ;
      RECT 0.680000 471.390000 538.390000 471.810000 ;
      RECT 0.000000 468.210000 538.390000 471.390000 ;
      RECT 0.680000 467.790000 538.390000 468.210000 ;
      RECT 0.000000 464.410000 538.390000 467.790000 ;
      RECT 0.680000 463.990000 538.390000 464.410000 ;
      RECT 0.000000 460.810000 538.390000 463.990000 ;
      RECT 0.680000 460.390000 538.390000 460.810000 ;
      RECT 0.000000 457.010000 538.390000 460.390000 ;
      RECT 0.680000 456.590000 538.390000 457.010000 ;
      RECT 0.000000 453.410000 538.390000 456.590000 ;
      RECT 0.680000 452.990000 538.390000 453.410000 ;
      RECT 0.000000 449.610000 538.390000 452.990000 ;
      RECT 0.680000 449.190000 538.390000 449.610000 ;
      RECT 0.000000 446.010000 538.390000 449.190000 ;
      RECT 0.680000 445.590000 538.390000 446.010000 ;
      RECT 0.000000 442.410000 538.390000 445.590000 ;
      RECT 0.680000 441.990000 538.390000 442.410000 ;
      RECT 0.000000 438.610000 538.390000 441.990000 ;
      RECT 0.680000 438.190000 538.390000 438.610000 ;
      RECT 0.000000 435.010000 538.390000 438.190000 ;
      RECT 0.680000 434.590000 538.390000 435.010000 ;
      RECT 0.000000 431.210000 538.390000 434.590000 ;
      RECT 0.680000 430.790000 538.390000 431.210000 ;
      RECT 0.000000 427.610000 538.390000 430.790000 ;
      RECT 0.680000 427.190000 538.390000 427.610000 ;
      RECT 0.000000 424.010000 538.390000 427.190000 ;
      RECT 0.680000 423.590000 538.390000 424.010000 ;
      RECT 0.000000 420.210000 538.390000 423.590000 ;
      RECT 0.680000 419.790000 538.390000 420.210000 ;
      RECT 0.000000 416.610000 538.390000 419.790000 ;
      RECT 0.680000 416.190000 538.390000 416.610000 ;
      RECT 0.000000 412.810000 538.390000 416.190000 ;
      RECT 0.680000 412.390000 538.390000 412.810000 ;
      RECT 0.000000 409.210000 538.390000 412.390000 ;
      RECT 0.680000 408.790000 538.390000 409.210000 ;
      RECT 0.000000 405.410000 538.390000 408.790000 ;
      RECT 0.680000 404.990000 538.390000 405.410000 ;
      RECT 0.000000 401.810000 538.390000 404.990000 ;
      RECT 0.680000 401.390000 538.390000 401.810000 ;
      RECT 0.000000 398.210000 538.390000 401.390000 ;
      RECT 0.680000 397.790000 538.390000 398.210000 ;
      RECT 0.000000 394.410000 538.390000 397.790000 ;
      RECT 0.680000 393.990000 538.390000 394.410000 ;
      RECT 0.000000 390.810000 538.390000 393.990000 ;
      RECT 0.680000 390.390000 538.390000 390.810000 ;
      RECT 0.000000 387.010000 538.390000 390.390000 ;
      RECT 0.680000 386.590000 538.390000 387.010000 ;
      RECT 0.000000 383.410000 538.390000 386.590000 ;
      RECT 0.680000 382.990000 538.390000 383.410000 ;
      RECT 0.000000 379.810000 538.390000 382.990000 ;
      RECT 0.680000 379.390000 538.390000 379.810000 ;
      RECT 0.000000 376.010000 538.390000 379.390000 ;
      RECT 0.680000 375.590000 538.390000 376.010000 ;
      RECT 0.000000 372.410000 538.390000 375.590000 ;
      RECT 0.680000 371.990000 538.390000 372.410000 ;
      RECT 0.000000 368.610000 538.390000 371.990000 ;
      RECT 0.680000 368.190000 538.390000 368.610000 ;
      RECT 0.000000 365.010000 538.390000 368.190000 ;
      RECT 0.680000 364.590000 538.390000 365.010000 ;
      RECT 0.000000 361.210000 538.390000 364.590000 ;
      RECT 0.680000 360.790000 538.390000 361.210000 ;
      RECT 0.000000 357.610000 538.390000 360.790000 ;
      RECT 0.680000 357.190000 538.390000 357.610000 ;
      RECT 0.000000 354.010000 538.390000 357.190000 ;
      RECT 0.680000 353.590000 538.390000 354.010000 ;
      RECT 0.000000 350.210000 538.390000 353.590000 ;
      RECT 0.680000 349.790000 538.390000 350.210000 ;
      RECT 0.000000 346.610000 538.390000 349.790000 ;
      RECT 0.680000 346.190000 538.390000 346.610000 ;
      RECT 0.000000 342.810000 538.390000 346.190000 ;
      RECT 0.680000 342.390000 538.390000 342.810000 ;
      RECT 0.000000 339.210000 538.390000 342.390000 ;
      RECT 0.680000 338.790000 538.390000 339.210000 ;
      RECT 0.000000 335.610000 538.390000 338.790000 ;
      RECT 0.680000 335.190000 538.390000 335.610000 ;
      RECT 0.000000 331.810000 538.390000 335.190000 ;
      RECT 0.680000 331.390000 538.390000 331.810000 ;
      RECT 0.000000 328.210000 538.390000 331.390000 ;
      RECT 0.680000 327.790000 538.390000 328.210000 ;
      RECT 0.000000 324.410000 538.390000 327.790000 ;
      RECT 0.680000 323.990000 538.390000 324.410000 ;
      RECT 0.000000 320.810000 538.390000 323.990000 ;
      RECT 0.680000 320.390000 538.390000 320.810000 ;
      RECT 0.000000 317.010000 538.390000 320.390000 ;
      RECT 0.680000 316.590000 538.390000 317.010000 ;
      RECT 0.000000 313.410000 538.390000 316.590000 ;
      RECT 0.680000 312.990000 538.390000 313.410000 ;
      RECT 0.000000 309.810000 538.390000 312.990000 ;
      RECT 0.680000 309.390000 538.390000 309.810000 ;
      RECT 0.000000 306.010000 538.390000 309.390000 ;
      RECT 0.680000 305.590000 538.390000 306.010000 ;
      RECT 0.000000 302.410000 538.390000 305.590000 ;
      RECT 0.680000 301.990000 538.390000 302.410000 ;
      RECT 0.000000 298.610000 538.390000 301.990000 ;
      RECT 0.680000 298.190000 538.390000 298.610000 ;
      RECT 0.000000 295.010000 538.390000 298.190000 ;
      RECT 0.680000 294.590000 538.390000 295.010000 ;
      RECT 0.000000 291.410000 538.390000 294.590000 ;
      RECT 0.680000 290.990000 538.390000 291.410000 ;
      RECT 0.000000 287.610000 538.390000 290.990000 ;
      RECT 0.680000 287.190000 538.390000 287.610000 ;
      RECT 0.000000 284.010000 538.390000 287.190000 ;
      RECT 0.680000 283.590000 538.390000 284.010000 ;
      RECT 0.000000 280.210000 538.390000 283.590000 ;
      RECT 0.680000 279.790000 538.390000 280.210000 ;
      RECT 0.000000 276.610000 538.390000 279.790000 ;
      RECT 0.680000 276.190000 538.390000 276.610000 ;
      RECT 0.000000 272.810000 538.390000 276.190000 ;
      RECT 0.680000 272.390000 538.390000 272.810000 ;
      RECT 0.000000 269.210000 538.390000 272.390000 ;
      RECT 0.680000 268.790000 538.390000 269.210000 ;
      RECT 0.000000 265.610000 538.390000 268.790000 ;
      RECT 0.680000 265.190000 538.390000 265.610000 ;
      RECT 0.000000 261.810000 538.390000 265.190000 ;
      RECT 0.680000 261.390000 538.390000 261.810000 ;
      RECT 0.000000 258.210000 538.390000 261.390000 ;
      RECT 0.680000 257.790000 538.390000 258.210000 ;
      RECT 0.000000 254.410000 538.390000 257.790000 ;
      RECT 0.680000 253.990000 538.390000 254.410000 ;
      RECT 0.000000 250.810000 538.390000 253.990000 ;
      RECT 0.680000 250.390000 538.390000 250.810000 ;
      RECT 0.000000 247.010000 538.390000 250.390000 ;
      RECT 0.680000 246.590000 538.390000 247.010000 ;
      RECT 0.000000 243.410000 538.390000 246.590000 ;
      RECT 0.680000 242.990000 538.390000 243.410000 ;
      RECT 0.000000 239.810000 538.390000 242.990000 ;
      RECT 0.680000 239.390000 538.390000 239.810000 ;
      RECT 0.000000 236.010000 538.390000 239.390000 ;
      RECT 0.680000 235.590000 538.390000 236.010000 ;
      RECT 0.000000 232.410000 538.390000 235.590000 ;
      RECT 0.680000 231.990000 538.390000 232.410000 ;
      RECT 0.000000 228.610000 538.390000 231.990000 ;
      RECT 0.680000 228.190000 538.390000 228.610000 ;
      RECT 0.000000 225.010000 538.390000 228.190000 ;
      RECT 0.680000 224.590000 538.390000 225.010000 ;
      RECT 0.000000 221.410000 538.390000 224.590000 ;
      RECT 0.680000 220.990000 538.390000 221.410000 ;
      RECT 0.000000 217.610000 538.390000 220.990000 ;
      RECT 0.680000 217.190000 538.390000 217.610000 ;
      RECT 0.000000 214.010000 538.390000 217.190000 ;
      RECT 0.680000 213.590000 538.390000 214.010000 ;
      RECT 0.000000 210.210000 538.390000 213.590000 ;
      RECT 0.680000 209.790000 538.390000 210.210000 ;
      RECT 0.000000 206.610000 538.390000 209.790000 ;
      RECT 0.680000 206.190000 538.390000 206.610000 ;
      RECT 0.000000 202.810000 538.390000 206.190000 ;
      RECT 0.680000 202.390000 538.390000 202.810000 ;
      RECT 0.000000 199.210000 538.390000 202.390000 ;
      RECT 0.680000 198.790000 538.390000 199.210000 ;
      RECT 0.000000 195.610000 538.390000 198.790000 ;
      RECT 0.680000 195.190000 538.390000 195.610000 ;
      RECT 0.000000 191.810000 538.390000 195.190000 ;
      RECT 0.680000 191.390000 538.390000 191.810000 ;
      RECT 0.000000 188.210000 538.390000 191.390000 ;
      RECT 0.680000 187.790000 538.390000 188.210000 ;
      RECT 0.000000 184.410000 538.390000 187.790000 ;
      RECT 0.680000 183.990000 538.390000 184.410000 ;
      RECT 0.000000 180.810000 538.390000 183.990000 ;
      RECT 0.680000 180.390000 538.390000 180.810000 ;
      RECT 0.000000 177.210000 538.390000 180.390000 ;
      RECT 0.680000 176.790000 538.390000 177.210000 ;
      RECT 0.000000 173.410000 538.390000 176.790000 ;
      RECT 0.680000 172.990000 538.390000 173.410000 ;
      RECT 0.000000 169.810000 538.390000 172.990000 ;
      RECT 0.680000 169.390000 538.390000 169.810000 ;
      RECT 0.000000 166.010000 538.390000 169.390000 ;
      RECT 0.680000 165.590000 538.390000 166.010000 ;
      RECT 0.000000 162.410000 538.390000 165.590000 ;
      RECT 0.680000 161.990000 538.390000 162.410000 ;
      RECT 0.000000 158.610000 538.390000 161.990000 ;
      RECT 0.680000 158.190000 538.390000 158.610000 ;
      RECT 0.000000 155.010000 538.390000 158.190000 ;
      RECT 0.680000 154.590000 538.390000 155.010000 ;
      RECT 0.000000 151.410000 538.390000 154.590000 ;
      RECT 0.680000 150.990000 538.390000 151.410000 ;
      RECT 0.000000 147.610000 538.390000 150.990000 ;
      RECT 0.680000 147.190000 538.390000 147.610000 ;
      RECT 0.000000 144.010000 538.390000 147.190000 ;
      RECT 0.680000 143.590000 538.390000 144.010000 ;
      RECT 0.000000 140.210000 538.390000 143.590000 ;
      RECT 0.680000 139.790000 538.390000 140.210000 ;
      RECT 0.000000 136.610000 538.390000 139.790000 ;
      RECT 0.680000 136.190000 538.390000 136.610000 ;
      RECT 0.000000 133.010000 538.390000 136.190000 ;
      RECT 0.680000 132.590000 538.390000 133.010000 ;
      RECT 0.000000 129.210000 538.390000 132.590000 ;
      RECT 0.680000 128.790000 538.390000 129.210000 ;
      RECT 0.000000 125.610000 538.390000 128.790000 ;
      RECT 0.680000 125.190000 538.390000 125.610000 ;
      RECT 0.000000 121.810000 538.390000 125.190000 ;
      RECT 0.680000 121.390000 538.390000 121.810000 ;
      RECT 0.000000 118.210000 538.390000 121.390000 ;
      RECT 0.680000 117.790000 538.390000 118.210000 ;
      RECT 0.000000 114.410000 538.390000 117.790000 ;
      RECT 0.680000 113.990000 538.390000 114.410000 ;
      RECT 0.000000 110.810000 538.390000 113.990000 ;
      RECT 0.680000 110.390000 538.390000 110.810000 ;
      RECT 0.000000 107.210000 538.390000 110.390000 ;
      RECT 0.680000 106.790000 538.390000 107.210000 ;
      RECT 0.000000 103.410000 538.390000 106.790000 ;
      RECT 0.680000 102.990000 538.390000 103.410000 ;
      RECT 0.000000 99.810000 538.390000 102.990000 ;
      RECT 0.680000 99.390000 538.390000 99.810000 ;
      RECT 0.000000 96.010000 538.390000 99.390000 ;
      RECT 0.680000 95.590000 538.390000 96.010000 ;
      RECT 0.000000 92.410000 538.390000 95.590000 ;
      RECT 0.680000 91.990000 538.390000 92.410000 ;
      RECT 0.000000 88.810000 538.390000 91.990000 ;
      RECT 0.680000 88.390000 538.390000 88.810000 ;
      RECT 0.000000 85.010000 538.390000 88.390000 ;
      RECT 0.680000 84.590000 538.390000 85.010000 ;
      RECT 0.000000 81.410000 538.390000 84.590000 ;
      RECT 0.680000 80.990000 538.390000 81.410000 ;
      RECT 0.000000 77.610000 538.390000 80.990000 ;
      RECT 0.680000 77.190000 538.390000 77.610000 ;
      RECT 0.000000 74.010000 538.390000 77.190000 ;
      RECT 0.680000 73.590000 538.390000 74.010000 ;
      RECT 0.000000 70.210000 538.390000 73.590000 ;
      RECT 0.680000 69.790000 538.390000 70.210000 ;
      RECT 0.000000 66.610000 538.390000 69.790000 ;
      RECT 0.680000 66.190000 538.390000 66.610000 ;
      RECT 0.000000 63.010000 538.390000 66.190000 ;
      RECT 0.680000 62.590000 538.390000 63.010000 ;
      RECT 0.000000 59.210000 538.390000 62.590000 ;
      RECT 0.680000 58.790000 538.390000 59.210000 ;
      RECT 0.000000 55.610000 538.390000 58.790000 ;
      RECT 0.680000 55.190000 538.390000 55.610000 ;
      RECT 0.000000 51.810000 538.390000 55.190000 ;
      RECT 0.680000 51.390000 538.390000 51.810000 ;
      RECT 0.000000 48.210000 538.390000 51.390000 ;
      RECT 0.680000 47.790000 538.390000 48.210000 ;
      RECT 0.000000 44.610000 538.390000 47.790000 ;
      RECT 0.680000 44.190000 538.390000 44.610000 ;
      RECT 0.000000 40.810000 538.390000 44.190000 ;
      RECT 0.680000 40.390000 538.390000 40.810000 ;
      RECT 0.000000 37.210000 538.390000 40.390000 ;
      RECT 0.680000 36.790000 538.390000 37.210000 ;
      RECT 0.000000 33.410000 538.390000 36.790000 ;
      RECT 0.680000 32.990000 538.390000 33.410000 ;
      RECT 0.000000 29.810000 538.390000 32.990000 ;
      RECT 0.680000 29.390000 538.390000 29.810000 ;
      RECT 0.000000 26.010000 538.390000 29.390000 ;
      RECT 0.680000 25.590000 538.390000 26.010000 ;
      RECT 0.000000 22.410000 538.390000 25.590000 ;
      RECT 0.680000 21.990000 538.390000 22.410000 ;
      RECT 0.000000 18.810000 538.390000 21.990000 ;
      RECT 0.680000 18.390000 538.390000 18.810000 ;
      RECT 0.000000 15.010000 538.390000 18.390000 ;
      RECT 0.680000 14.590000 538.390000 15.010000 ;
      RECT 0.000000 11.410000 538.390000 14.590000 ;
      RECT 0.680000 10.990000 538.390000 11.410000 ;
      RECT 0.000000 7.610000 538.390000 10.990000 ;
      RECT 0.680000 7.190000 538.390000 7.610000 ;
      RECT 0.000000 4.010000 538.390000 7.190000 ;
      RECT 0.680000 3.590000 538.390000 4.010000 ;
      RECT 0.000000 0.640000 538.390000 3.590000 ;
      RECT 0.000000 0.410000 0.550000 0.640000 ;
      RECT 535.250000 0.000000 538.150000 0.640000 ;
      RECT 531.850000 0.000000 534.950000 0.640000 ;
      RECT 528.450000 0.000000 531.550000 0.640000 ;
      RECT 525.050000 0.000000 528.150000 0.640000 ;
      RECT 521.650000 0.000000 524.750000 0.640000 ;
      RECT 518.250000 0.000000 521.350000 0.640000 ;
      RECT 514.850000 0.000000 517.950000 0.640000 ;
      RECT 511.450000 0.000000 514.550000 0.640000 ;
      RECT 508.050000 0.000000 511.150000 0.640000 ;
      RECT 504.650000 0.000000 507.750000 0.640000 ;
      RECT 501.250000 0.000000 504.350000 0.640000 ;
      RECT 497.850000 0.000000 500.950000 0.640000 ;
      RECT 494.450000 0.000000 497.550000 0.640000 ;
      RECT 491.250000 0.000000 494.150000 0.640000 ;
      RECT 487.850000 0.000000 490.950000 0.640000 ;
      RECT 484.450000 0.000000 487.550000 0.640000 ;
      RECT 481.050000 0.000000 484.150000 0.640000 ;
      RECT 477.650000 0.000000 480.750000 0.640000 ;
      RECT 474.250000 0.000000 477.350000 0.640000 ;
      RECT 470.850000 0.000000 473.950000 0.640000 ;
      RECT 467.450000 0.000000 470.550000 0.640000 ;
      RECT 464.050000 0.000000 467.150000 0.640000 ;
      RECT 460.650000 0.000000 463.750000 0.640000 ;
      RECT 457.250000 0.000000 460.350000 0.640000 ;
      RECT 453.850000 0.000000 456.950000 0.640000 ;
      RECT 450.450000 0.000000 453.550000 0.640000 ;
      RECT 447.250000 0.000000 450.150000 0.640000 ;
      RECT 443.850000 0.000000 446.950000 0.640000 ;
      RECT 440.450000 0.000000 443.550000 0.640000 ;
      RECT 437.050000 0.000000 440.150000 0.640000 ;
      RECT 433.650000 0.000000 436.750000 0.640000 ;
      RECT 430.250000 0.000000 433.350000 0.640000 ;
      RECT 426.850000 0.000000 429.950000 0.640000 ;
      RECT 423.450000 0.000000 426.550000 0.640000 ;
      RECT 420.050000 0.000000 423.150000 0.640000 ;
      RECT 416.650000 0.000000 419.750000 0.640000 ;
      RECT 413.250000 0.000000 416.350000 0.640000 ;
      RECT 409.850000 0.000000 412.950000 0.640000 ;
      RECT 406.450000 0.000000 409.550000 0.640000 ;
      RECT 403.250000 0.000000 406.150000 0.640000 ;
      RECT 399.850000 0.000000 402.950000 0.640000 ;
      RECT 396.450000 0.000000 399.550000 0.640000 ;
      RECT 393.050000 0.000000 396.150000 0.640000 ;
      RECT 389.650000 0.000000 392.750000 0.640000 ;
      RECT 386.250000 0.000000 389.350000 0.640000 ;
      RECT 382.850000 0.000000 385.950000 0.640000 ;
      RECT 379.450000 0.000000 382.550000 0.640000 ;
      RECT 376.050000 0.000000 379.150000 0.640000 ;
      RECT 372.650000 0.000000 375.750000 0.640000 ;
      RECT 369.250000 0.000000 372.350000 0.640000 ;
      RECT 365.850000 0.000000 368.950000 0.640000 ;
      RECT 362.450000 0.000000 365.550000 0.640000 ;
      RECT 359.250000 0.000000 362.150000 0.640000 ;
      RECT 355.850000 0.000000 358.950000 0.640000 ;
      RECT 352.450000 0.000000 355.550000 0.640000 ;
      RECT 349.050000 0.000000 352.150000 0.640000 ;
      RECT 345.650000 0.000000 348.750000 0.640000 ;
      RECT 342.250000 0.000000 345.350000 0.640000 ;
      RECT 338.850000 0.000000 341.950000 0.640000 ;
      RECT 335.450000 0.000000 338.550000 0.640000 ;
      RECT 332.050000 0.000000 335.150000 0.640000 ;
      RECT 328.650000 0.000000 331.750000 0.640000 ;
      RECT 325.250000 0.000000 328.350000 0.640000 ;
      RECT 321.850000 0.000000 324.950000 0.640000 ;
      RECT 318.450000 0.000000 321.550000 0.640000 ;
      RECT 315.050000 0.000000 318.150000 0.640000 ;
      RECT 311.850000 0.000000 314.750000 0.640000 ;
      RECT 308.450000 0.000000 311.550000 0.640000 ;
      RECT 305.050000 0.000000 308.150000 0.640000 ;
      RECT 301.650000 0.000000 304.750000 0.640000 ;
      RECT 298.250000 0.000000 301.350000 0.640000 ;
      RECT 294.850000 0.000000 297.950000 0.640000 ;
      RECT 291.450000 0.000000 294.550000 0.640000 ;
      RECT 288.050000 0.000000 291.150000 0.640000 ;
      RECT 284.650000 0.000000 287.750000 0.640000 ;
      RECT 281.250000 0.000000 284.350000 0.640000 ;
      RECT 277.850000 0.000000 280.950000 0.640000 ;
      RECT 274.450000 0.000000 277.550000 0.640000 ;
      RECT 271.050000 0.000000 274.150000 0.640000 ;
      RECT 267.850000 0.000000 270.750000 0.640000 ;
      RECT 264.450000 0.000000 267.550000 0.640000 ;
      RECT 261.050000 0.000000 264.150000 0.640000 ;
      RECT 257.650000 0.000000 260.750000 0.640000 ;
      RECT 254.250000 0.000000 257.350000 0.640000 ;
      RECT 250.850000 0.000000 253.950000 0.640000 ;
      RECT 247.450000 0.000000 250.550000 0.640000 ;
      RECT 244.050000 0.000000 247.150000 0.640000 ;
      RECT 240.650000 0.000000 243.750000 0.640000 ;
      RECT 237.250000 0.000000 240.350000 0.640000 ;
      RECT 233.850000 0.000000 236.950000 0.640000 ;
      RECT 230.450000 0.000000 233.550000 0.640000 ;
      RECT 227.050000 0.000000 230.150000 0.640000 ;
      RECT 223.850000 0.000000 226.750000 0.640000 ;
      RECT 220.450000 0.000000 223.550000 0.640000 ;
      RECT 217.050000 0.000000 220.150000 0.640000 ;
      RECT 213.650000 0.000000 216.750000 0.640000 ;
      RECT 210.250000 0.000000 213.350000 0.640000 ;
      RECT 206.850000 0.000000 209.950000 0.640000 ;
      RECT 203.450000 0.000000 206.550000 0.640000 ;
      RECT 200.050000 0.000000 203.150000 0.640000 ;
      RECT 196.650000 0.000000 199.750000 0.640000 ;
      RECT 193.250000 0.000000 196.350000 0.640000 ;
      RECT 189.850000 0.000000 192.950000 0.640000 ;
      RECT 186.450000 0.000000 189.550000 0.640000 ;
      RECT 183.050000 0.000000 186.150000 0.640000 ;
      RECT 179.850000 0.000000 182.750000 0.640000 ;
      RECT 176.450000 0.000000 179.550000 0.640000 ;
      RECT 173.050000 0.000000 176.150000 0.640000 ;
      RECT 169.650000 0.000000 172.750000 0.640000 ;
      RECT 166.250000 0.000000 169.350000 0.640000 ;
      RECT 162.850000 0.000000 165.950000 0.640000 ;
      RECT 159.450000 0.000000 162.550000 0.640000 ;
      RECT 156.050000 0.000000 159.150000 0.640000 ;
      RECT 152.650000 0.000000 155.750000 0.640000 ;
      RECT 149.250000 0.000000 152.350000 0.640000 ;
      RECT 145.850000 0.000000 148.950000 0.640000 ;
      RECT 142.450000 0.000000 145.550000 0.640000 ;
      RECT 139.050000 0.000000 142.150000 0.640000 ;
      RECT 135.650000 0.000000 138.750000 0.640000 ;
      RECT 132.450000 0.000000 135.350000 0.640000 ;
      RECT 129.050000 0.000000 132.150000 0.640000 ;
      RECT 125.650000 0.000000 128.750000 0.640000 ;
      RECT 122.250000 0.000000 125.350000 0.640000 ;
      RECT 118.850000 0.000000 121.950000 0.640000 ;
      RECT 115.450000 0.000000 118.550000 0.640000 ;
      RECT 112.050000 0.000000 115.150000 0.640000 ;
      RECT 108.650000 0.000000 111.750000 0.640000 ;
      RECT 105.250000 0.000000 108.350000 0.640000 ;
      RECT 101.850000 0.000000 104.950000 0.640000 ;
      RECT 98.450000 0.000000 101.550000 0.640000 ;
      RECT 95.050000 0.000000 98.150000 0.640000 ;
      RECT 91.650000 0.000000 94.750000 0.640000 ;
      RECT 88.450000 0.000000 91.350000 0.640000 ;
      RECT 85.050000 0.000000 88.150000 0.640000 ;
      RECT 81.650000 0.000000 84.750000 0.640000 ;
      RECT 78.250000 0.000000 81.350000 0.640000 ;
      RECT 74.850000 0.000000 77.950000 0.640000 ;
      RECT 71.450000 0.000000 74.550000 0.640000 ;
      RECT 68.050000 0.000000 71.150000 0.640000 ;
      RECT 64.650000 0.000000 67.750000 0.640000 ;
      RECT 61.250000 0.000000 64.350000 0.640000 ;
      RECT 57.850000 0.000000 60.950000 0.640000 ;
      RECT 54.450000 0.000000 57.550000 0.640000 ;
      RECT 51.050000 0.000000 54.150000 0.640000 ;
      RECT 47.650000 0.000000 50.750000 0.640000 ;
      RECT 44.450000 0.000000 47.350000 0.640000 ;
      RECT 41.050000 0.000000 44.150000 0.640000 ;
      RECT 37.650000 0.000000 40.750000 0.640000 ;
      RECT 34.250000 0.000000 37.350000 0.640000 ;
      RECT 30.850000 0.000000 33.950000 0.640000 ;
      RECT 27.450000 0.000000 30.550000 0.640000 ;
      RECT 24.050000 0.000000 27.150000 0.640000 ;
      RECT 20.650000 0.000000 23.750000 0.640000 ;
      RECT 17.250000 0.000000 20.350000 0.640000 ;
      RECT 13.850000 0.000000 16.950000 0.640000 ;
      RECT 10.450000 0.000000 13.550000 0.640000 ;
      RECT 7.050000 0.000000 10.150000 0.640000 ;
      RECT 3.650000 0.000000 6.750000 0.640000 ;
      RECT 0.850000 0.000000 3.350000 0.640000 ;
    LAYER M5 ;
      RECT 0.000000 0.000000 538.390000 538.200000 ;
    LAYER M6 ;
      RECT 0.000000 0.000000 538.390000 538.200000 ;
    LAYER M7 ;
      RECT 0.000000 0.000000 538.390000 538.200000 ;
    LAYER M8 ;
      RECT 0.000000 0.000000 538.390000 538.200000 ;
  END
END fullchip

END LIBRARY
