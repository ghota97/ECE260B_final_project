/home/linux/ieng6/ee260bwi22/public/PDKdata/lef/tcbn65gplus_8lmT2.lef